interface dec_intf;
logic [2:0]i;
logic [7:0]d;
endinterface
