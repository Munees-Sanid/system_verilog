interface dff_if;
logic clk,rst;
logic d; // input of d flip flop
logic q; // output of d flip flop
  
endinterface
