interface dff_if;
logic clk,rst;
logic din;
logic dout;
  
endinterface
