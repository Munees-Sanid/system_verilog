module tb;
logic a;
bit b;
byte c;
longint d;
int e;
shortint f;
initial begin 
$display("default value of logic is %b",$bits)
