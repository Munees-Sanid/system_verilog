module tb;
int a;
real b;
initial begin
$display($bits(a));
$display($bits(b));
end
endmodule
