interface tff_if;
logic clk,rst;
logic t; // input of t flip flop
logic q; // output of t flip flop
  
endinterface
