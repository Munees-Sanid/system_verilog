interface enc_intf;
logic [7:0]i;
logic [2:0]y;
endinterface
