interface comp_intf;
logic a,b;
logic eq,gt,lt;
endinterface
